----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12/26/2021 01:04:07 PM
-- Design Name: 
-- Module Name: keypad - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity KEYPAD is

GENERIC(
			FREQ_CLK : INTEGER := 125000000         --FRECUENCIA DE LA TARJETA
);


PORT(
	CLK 		  : IN  STD_LOGIC; 				   --RELOJ FPGA
	COLUMNAS   : IN  STD_LOGIC_VECTOR(3  DOWNTO 0); --PUERTO CONECTADO A LAS COLUMNAS DEL TECLADO
	FILAS 	  : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);  --PUERTO CONECTADO A LA FILAS DEL TECLADO
	BOTON_PRES : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); --PUERTO QUE INDICA LA TECLA QUE SE PRESION�"
	IND		  : OUT STD_LOGIC					   --BANDERA QUE INDICA CUANDO SE PRESION�" UNA TECLA (S�"LO DURA UN CICLO DE RELOJ)
);

end KEYPAD;

architecture Behavioral of KEYPAD is

CONSTANT DELAY_1MS  : INTEGER := (FREQ_CLK/1000)-1;
CONSTANT DELAY_10MS : INTEGER := (FREQ_CLK/100)-1;

SIGNAL CONTA_1MS 	: INTEGER RANGE 0 TO DELAY_1MS := 0;
SIGNAL BANDERA 	: STD_LOGIC := '0';
SIGNAL CONTA_10MS : INTEGER RANGE 0 TO DELAY_10MS := 0;
SIGNAL BANDERA2 	: STD_LOGIC := '0';

SIGNAL REG_B1  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B2  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B3  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B4  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B5  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B6  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B7  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B8  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B9  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B0  : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_BAS : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_BGA : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_A : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_B : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_C : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');
SIGNAL REG_D : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS=>'0');

SIGNAL FILA_REG_S : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS=>'0');
SIGNAL FILA : INTEGER RANGE 0 TO 3 := 0;

SIGNAL IND_S : STD_LOGIC := '0';
SIGNAL EDO : INTEGER RANGE 0 TO 1 := 0;

begin

FILAS <= FILA_REG_S;

--RETARDO 1 MS--
PROCESS(CLK)
BEGIN
IF RISING_EDGE(CLK) THEN
	CONTA_1MS <= CONTA_1MS+1;
	BANDERA <= '0';
	IF CONTA_1MS = DELAY_1MS THEN
		CONTA_1MS <= 0;
		BANDERA <= '1';
	END IF;
END IF;
END PROCESS;
----------------

--RETARDO 10 MS--
PROCESS(CLK)
BEGIN
IF RISING_EDGE(CLK) THEN
	CONTA_10MS <= CONTA_10MS+1;
	BANDERA2 <= '0';
	IF CONTA_10MS = DELAY_10MS THEN
		CONTA_10MS <= 0;
		BANDERA2 <= '1';
	END IF;
END IF;
END PROCESS;
----------------

--PROCESO QUE ACTIVA/BARRIDO CADA FILA CADA 10ms--
PROCESS(CLK, BANDERA2)
BEGIN
	IF RISING_EDGE(CLK) AND BANDERA2 = '1' THEN
		FILA <= FILA+1;
		IF FILA = 3 THEN
			FILA <= 0;
		END IF;
	END IF;
END PROCESS;

WITH FILA SELECT
	FILA_REG_S <= "1000" WHEN 0,
					  "0100" WHEN 1,
					  "0010" WHEN 2,
					  "0001" WHEN OTHERS;
-------------------------------				

----------PROCESO QUE EVITA EL EFECTO REBOTE DE LAS TECLAS----------------
--LLENA LOS REGISTROS CON '1' DEPENDIENDO EL BOT�"N QUE SE HAYA PRESIONADO--
PROCESS(CLK,BANDERA)
BEGIN
	IF RISING_EDGE(CLK) AND BANDERA = '1' THEN
	    IF COLUMNAS = "0000" THEN
	          REG_B1 <= (others => '0');
	          REG_B2 <= (others => '0');
	          REG_B3 <= (others => '0');
	          REG_B4 <= (others => '0');
	          REG_B5 <= (others => '0');
	          REG_B6 <= (others => '0');
	          REG_B7 <= (others => '0');
	          REG_B8 <= (others => '0');
	          REG_B9 <= (others => '0');
	          REG_B0 <= (others => '0');
	          REG_A <= (others => '0');
	          REG_B <= (others => '0');
	          REG_C <= (others => '0');
	          REG_D <= (others => '0');
	          REG_BGA <= (others => '0');
	          REG_BAS <= (others => '0');
		ELSIF FILA_REG_S = "1000" THEN --PRIMERA FILA DE BOTONES
			REG_B1 <= REG_B1(6 DOWNTO 0)&COLUMNAS(3);
			REG_B2 <= REG_B2(6 DOWNTO 0)&COLUMNAS(2);
			REG_B3 <= REG_B3(6 DOWNTO 0)&COLUMNAS(1);
			REG_A <= REG_A(6 DOWNTO 0)&COLUMNAS(0);
		ELSIF FILA_REG_S = "0100" THEN --SEGUNDA FILA DE BOTONES
			REG_B4 <= REG_B4(6 DOWNTO 0)&COLUMNAS(3);
			REG_B5 <= REG_B5(6 DOWNTO 0)&COLUMNAS(2);
			REG_B6 <= REG_B6(6 DOWNTO 0)&COLUMNAS(1);
			REG_B <= REG_B(6 DOWNTO 0)&COLUMNAS(0);
		ELSIF FILA_REG_S = "0010" THEN --TERCERA FILA DE BOTONES
			REG_B7 <= REG_B7(6 DOWNTO 0)&COLUMNAS(3);
			REG_B8 <= REG_B8(6 DOWNTO 0)&COLUMNAS(2);
			REG_B9 <= REG_B9(6 DOWNTO 0)&COLUMNAS(1);
		    REG_C <= REG_C(6 DOWNTO 0)&COLUMNAS(0);
		ELSIF FILA_REG_S = "0001" THEN --CUARTA FILA DE BOTONES
			REG_BAS <= REG_BAS(6 DOWNTO 0)&COLUMNAS(3);
			REG_B0  <= REG_B0(6 DOWNTO 0)&COLUMNAS(2);
			REG_BGA <= REG_BGA(6 DOWNTO 0)&COLUMNAS(1);
			  REG_D <= REG_D(6 DOWNTO 0)&COLUMNAS(0);
		END IF;
	END IF;
END PROCESS;
----------------------------------------------------------------------------

--MANDA EL DATO A LA SALIDA--
PROCESS(CLK)
BEGIN
	IF RISING_EDGE(CLK) THEN
		IF 	REG_B0  	= "11111111" THEN BOTON_PRES <= X"30"; IND_S <= '1';
		ELSIF REG_B1 	= "11111111" THEN BOTON_PRES <= X"31"; IND_S <= '1';
		ELSIF	REG_B2 	= "11111111" THEN BOTON_PRES <= X"32"; IND_S <= '1';
		ELSIF	REG_B3 	= "11111111" THEN BOTON_PRES <= X"33"; IND_S <= '1';
		ELSIF	REG_B4 	= "11111111" THEN BOTON_PRES <= X"34"; IND_S <= '1';
		ELSIF	REG_B5 	= "11111111" THEN BOTON_PRES <= X"35"; IND_S <= '1';
		ELSIF	REG_B6 	= "11111111" THEN BOTON_PRES <= X"36"; IND_S <= '1';
		ELSIF	REG_B7 	= "11111111" THEN BOTON_PRES <= X"37"; IND_S <= '1';
		ELSIF	REG_B8 	= "11111111" THEN BOTON_PRES <= X"38"; IND_S <= '1';
		ELSIF	REG_B9 	= "11111111" THEN BOTON_PRES <= X"39"; IND_S <= '1';
		ELSIF	REG_A 	= "11111111" THEN BOTON_PRES <= X"41"; IND_S <= '1';
		ELSIF	REG_B 	= "11111111" THEN BOTON_PRES <= X"42"; IND_S <= '1';
		ELSIF	REG_C 	= "11111111" THEN BOTON_PRES <= X"43"; IND_S <= '1';
		ELSIF	REG_D 	= "11111111" THEN BOTON_PRES <= X"44"; IND_S <= '1'; 
		ELSIF	REG_BAS 	= "11111111" THEN BOTON_PRES <= X"2A"; IND_S <= '1';
		ELSIF	REG_BGA 	= "11111111" THEN BOTON_PRES <= X"23"; IND_S <= '1';
		ELSE IND_S <= '0';
		END IF;
	END IF;
END PROCESS;
-----------------------------

--M�?QUINA DE ESTADOS PARA LA BANDERA--
PROCESS(IND_S,CLK)
BEGIN
	IF RISING_EDGE(CLK) THEN
				IND <= IND_S;
    END IF;
END PROCESS;
--------------------------------------


end Behavioral;